`ifndef TEST_UTILS_PARAMS
`define TEST_UTILS_PARAMS

//------------------------------------------------------------------------
// Console colors
//------------------------------------------------------------------------

`define CLI_RED    "\033[31m"
`define CLI_GREEN  "\033[32m"
`define CLI_YELLOW "\033[33m"
`define CLI_BLUE   "\033[34m"
`define CLI_RESET  "\033[0m"

//------------------------------------------------------------------------
// Common values
//------------------------------------------------------------------------
`define TB_CASE_DRAIN_TIME 100

`endif
